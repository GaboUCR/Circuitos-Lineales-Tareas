C:\Users\gabri\Dropbox\University\Circuitos lineales 1\tareas\Tarea4\Simulaciones\circuit2.cir DC Analysis
* Converted From Micro Cap Source file to SPICE3
*
.FUNC DPWR(D) {I(D)*V(D)}
.FUNC BPWR(Q) {IC(Q)*VCE(Q)+IB(Q)*VBE(Q)}
.FUNC FPWR(M) {ID(M)*VDS(M)}
.FUNC HOTD(D,MAX) {IF((V(D)*I(D)>MAX),1,0)}
.FUNC HOTB(Q,MAX) {IF((VCE(Q)*IC(Q)+IB(Q)*VBE(Q)>MAX),1,0)}
.FUNC HOTF(M,MAX) {IF((VDS(M)*ID(M)>MAX),1,0)}
.PARAM LOW3MIN={IMPORT(LOW3MIN.OUT,LOW3THRES)}
.PARAM HIGH3MAX={IMPORT(HIGH3MAX.OUT,HIGH3THRES)}
.PARAM LOWLVDS={IMPORT(LOWLVDS.OUT,LOWLIMIT)}
.PARAM HILVDS={IMPORT(HILVDS.OUT,HILIMIT)}
.PARAM LIMTLVDS={IMPORT(LIMTLVDS.OUT,LVDSLIMITS)}
.FUNC SKINAC(DCRES,RESISTIVITY,RELPERM,RADIUS) {((PI*RADIUS*RADIUS)/((PI*RADIUS*RADIUS)-PI*(RADIUS-SKINDEPTHAC(RESISTIVITY,RELPERM))**2))*DCRES}
.FUNC SKINDEPTHAC(RESISTIVITY,RELPERM) {503.3*(SQRT(RESISTIVITY/(RELPERM*F)))}
.FUNC SKINTR(DCRES,RESISTIVITY,RELPERM,RADIUS,FREQ) {((PI*RADIUS*RADIUS)/((PI*RADIUS*RADIUS)-PI*(RADIUS-SKINDEPTHTR(RESISTIVITY,RELPERM,FREQ))**2))*DCRES}
.FUNC SKINDEPTHTR(RESISTIVITY,RELPERM,FREQ) {503.3*(SQRT(RESISTIVITY/(RELPERM*FREQ)))}
E1 21 9 14 11 2
F1 4 6 VF1 1.2
G1 12 13 14 11 0.1
H1 15 17 VH1 {6}
I1 16 23 DC 0.5 
R1 0 1 30000
R2 2 0 30000
R3 3 0 10000
R4 4 1 20000
R5 3 4 10000
R7 4 2 30000
R8 1 4 10000
R9 3 5 20000
R10 6 5 30000
R11 4 6 10000
R12 4 9 20000
R13 2 9 10000
R14 2 9 20000
R15 3 5 20000
R16 9 5 10000
R17 10 5 10000
R18 5 11 30000
R19 12 11 10000
R20 15 13 30000
R21 16 13 10000
R22 15 10 20000
R23 17 10 20000
R24 19 17 30000
R25 19 16 10000
R26 20 19 20000
R27 21 20 10000
R28 2 9 30000
R29 2 16 20000
R30 8 16 10000
R31 2 8 20000
R32 8 16 30000
R33 18 16 20000
R34 8 22 10000
R35 22 23 30000
R36 22 23 20000
R37 22 24 30000
R38 16 23 20000
R39 25 24 20000
R40 24 26 30000
R41 23 25 10000
R42 25 27 10000
R43 27 28 10000
R44 27 12 20000
R45 26 14 10000
R46 28 14 30000
R47 14 11 20000
R48 12 11 30000
RE1 14 11 1G;added by E1
RG1 14 11 1G ;added by G1
V1 16 20 DC 20 
VF1 7 8 0 ;added by F1
VH1 18 7 0 ;added by H1
*
.LIB "C:\MC12\library\NOM.LIB"
*
*
.DC 0 0 0 0
*
.PROBE
.END
;$SpiceType=SPICE3
